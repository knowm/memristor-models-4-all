* Voltage Sources
V1 1 0 SIN(0V 0.5V 100Hz)

* Memristors
YMEMRISTOR mr1 1 0 mrm1 R_init=500

.MODEL mrm1 memristor (level=5 Roff=1500 Ron=500 Voff=0.27 Von=0.27 TAU=0.0001 PHI=0.8 SFA=0.0008 SFB=4 SRA=0.0008 SRB=4)

* Analysis Command
.TRAN .1ms .04s
* Output
.PRINT TRAN V(1) I(V1) N(YMEMRISTOR!mr1:R)

.END