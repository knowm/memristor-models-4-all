* test hys.va in DC, TRAN and Homotopy

V1 1 0 1 sin(0 0.7 1k)
Yhys H1 0 1

* DC analysis
.dc V1 -1 1 0.01
.print dc V(1) I(V1) N(Yhys!H1_ns)


* transient simulation
*.tran 1u 2m
*.print tran V(1) I(V1) N(Yhys!H1_ns)


