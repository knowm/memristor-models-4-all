
* Voltage Sources
V1 1 0 SIN(0V .25V 100Hz)

* Memristors
YMSSMEMRISTOR M1 1 0 

* Analysis Command
.TRAN .01ms 10ms
* Output
.PRINT TRAN V(1) I(V1) 


.END
